// A pro module for a comparator

module Comparator(

);

endmodule 